library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.Gates.all;

entity superscalar is
	port();
end entity;

architecture struct of superscalar is
begin

end architecture struct;