library IEEE;
use IEEE.std_logic_1164.all;

entity register_file is
	port ();
end entity register_file;

architecture trivial of register_file is
	begin
		

end architecture trivial;