library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.Gates.all;

entity rob is
    port(dispatch_word1, dispatch_word2: in std_logic_vector(len_PC +  downto 0); --I am assuming that each PC is
    );
end entity;
